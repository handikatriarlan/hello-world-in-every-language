// This is hello world verilog program.

module hello_world;

  initial begin
    $display("Hello, World!\n");
    $finish;
  end

endmodule
