module main

fn main() {
    println('Hello, World!')
}

# Execute this command to run the code : v run hello_world.v
